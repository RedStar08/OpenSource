library verilog;
use verilog.vl_types.all;
entity mux4_1tb is
end mux4_1tb;
