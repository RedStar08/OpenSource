library verilog;
use verilog.vl_types.all;
entity \_74LS138_tb\ is
end \_74LS138_tb\;
