module 74LS138_tb;
reg a;
reg b;
reg c;
wire [15:0]out;
	my4_16 my4_160(
		.a(a),
		.b(b),
		.c(c),
		.out(out)
	);
	
	initial begin
		a=0;b=0;c=0;d=0;
		#200;
		a=0;b=0;c=0;d=1;
		#200;
		a=0;b=0;c=1;d=0;
		#200;
		a=0;b=0;c=1;d=1;
		#200;
		
		a=0;b=1;c=0;d=0;
		#200;
		a=0;b=1;c=0;d=1;
		#200;
		a=0;b=1;c=1;d=0;
		#200;
		a=0;b=1;c=1;d=1;
		#200;
		
		a=1;b=0;c=0;d=0;
		#200;
		a=1;b=0;c=0;d=1;
		#200;
		a=1;b=0;c=1;d=0;
		#200;
		a=1;b=0;c=1;d=1;
		#200;
		
		a=1;b=1;c=0;d=0;
		#200;
		a=1;b=1;c=0;d=1;
		#200;
		a=1;b=1;c=1;d=0;
		#200;
		a=1;b=1;c=1;d=1;
		#200;
		
		$stop;	
	end
